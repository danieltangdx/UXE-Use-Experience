// xc_work/v/13.sv
// counter.v:0
// NOTE: This file corresponds to a module in the Hardware/DUT partition
`timescale 1ps/100fs
module _ixc_isc;
endmodule

