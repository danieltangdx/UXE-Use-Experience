library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity axis_delay is
  port (
    z : out std_logic ;
  a : in std_logic ) ;
end axis_delay ;
