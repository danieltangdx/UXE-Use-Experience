library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ixc_2xbuf is
  port (
    cout : out std_logic ;
  cin : in std_logic ) ;
end ixc_2xbuf ;
