library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity axis_busreg is
  port (
    z : inout std_logic ;
  DUMMY0 : inout std_logic ) ;
end axis_busreg ;
