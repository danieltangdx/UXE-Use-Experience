architecture module of ixc_bind is

begin
end module;
