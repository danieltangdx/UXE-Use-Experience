library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity IXC_MC_GSFIFO is
end IXC_MC_GSFIFO ;
