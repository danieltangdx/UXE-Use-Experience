library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ixc_osf_evcap is
  port (
    pvec : in std_logic ;
  pvecEv : out std_logic ) ;
  -- quickturn keep_net pvecEv
end ixc_osf_evcap ;
