library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ixc_asgn_cov_rst_pulse is
  port (
  rstsig : out std_logic ) ;
end ixc_asgn_cov_rst_pulse ;
