architecture module of IXC_ISF is

begin
end module;
