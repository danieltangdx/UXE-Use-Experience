library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity xc_top is
  generic (
    IXC_TIME : integer := 0
  ) ;
end xc_top ;
