// xc_work/v/7.sv
// /tools/cadence/UXE171_p98/tools.lnx86/etc/ixcom/IXCSF.sv:320
// NOTE: This file corresponds to a module in the Hardware/DUT partition
`timescale 1ps/100fs
module IXC_ISF;
endmodule

