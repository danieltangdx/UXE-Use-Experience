library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ixc_1xbufsrc is
  port (
    cout : out std_logic ;
  cin : in std_logic ) ;
end ixc_1xbufsrc ;
