
module xc_top ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire fclk;
wire _ET3_COMPILER_RESERVED_NAME_DUTPI_APPLY_;
wire _ET3_COMPILER_RESERVED_NAME_LBRKER_ON_;
wire callEmuPI;
wire [63:0] evalStepPI;
wire ckgHoldPI;
wire tbcHoldPI;
wire noOutputPI;
wire stopEmuPI;
wire oneStepPI;
wire stop1;
wire stop2;
wire stop4;
wire asyncCall;
wire isfWait;
wire osfWait;
wire sdlStop;
wire cpfStop;
wire eClk;
wire rClk;
wire bWait;
wire poBusy;
wire APPLY_PI;
wire lbrOnAll;
wire eClkv;
wire intr;
wire _zz_xmr0;
wire memWriteCmd;
wire dummyW;
wire _ET3_COMPILER_RESERVED_NAME_ORION_INTERRUPT_;
wire _ET3_COMPILER_RESERVED_NAME_DBI_APPLY_;
wire hotSwapOnPI;
wire sendPO;
wire tbcPO;
wire stop1PO;
wire stop2PO;
wire stop4PO;
wire stop3PO;
wire it_newBufPO;
wire stopSDLPO;
wire stopEmuPO;
wire stopCPFPO;
wire [63:0] remStepPO;
wire stop3;
wire stopSDL;
wire sdlEnable;
wire sdlHaltHwClk;
wire hwClkDbg;
wire hwClkDbgTime;
wire hwClkEnable;
wire hssReset;
wire tbcEnable;
wire [7:0] fclkPerEval;
wire evalOn;
wire evalOnOrig;
wire callEmuR;
wire eClkR;
wire callEmu;
wire callEmuD;
wire [63:0] eCount;
wire [63:0] evfCount;
wire [7:0] evalOnDExt;
wire [7:0] evalOnDCtl;
wire gfifoOff;
wire [63:0] simTime;
wire applyPiR;
wire dbiEvent;
wire FvUseOnly;
wire FvUseOnlyR;
wire eventOn;
wire mpSampleOv;
wire [7:0] poDelay;
wire lbrOn;
wire lbrOnD;
wire _zzmemWriteCmd;
wire dummyR;
supply0 n115;
supply1 n119;
supply0 n120;
supply1 n121;
supply1 n259;
Q_BUF U0 ( .A(n259), .Z(_ET3_COMPILER_RESERVED_NAME_DUTPI_APPLY_));
Q_BUF U1 ( .A(n115), .Z(it_newBufPO));
Q_BUF U2 ( .A(eventOn), .Z(mpSampleOv));
Q_BUF U3 ( .A(eCount[0]), .Z(remStepPO[0]));
Q_BUF U4 ( .A(eCount[1]), .Z(remStepPO[1]));
Q_BUF U5 ( .A(eCount[2]), .Z(remStepPO[2]));
Q_BUF U6 ( .A(eCount[3]), .Z(remStepPO[3]));
Q_BUF U7 ( .A(eCount[4]), .Z(remStepPO[4]));
Q_BUF U8 ( .A(eCount[5]), .Z(remStepPO[5]));
Q_BUF U9 ( .A(eCount[6]), .Z(remStepPO[6]));
Q_BUF U10 ( .A(eCount[7]), .Z(remStepPO[7]));
Q_BUF U11 ( .A(eCount[8]), .Z(remStepPO[8]));
Q_BUF U12 ( .A(eCount[9]), .Z(remStepPO[9]));
Q_BUF U13 ( .A(eCount[10]), .Z(remStepPO[10]));
Q_BUF U14 ( .A(eCount[11]), .Z(remStepPO[11]));
Q_BUF U15 ( .A(eCount[12]), .Z(remStepPO[12]));
Q_BUF U16 ( .A(eCount[13]), .Z(remStepPO[13]));
Q_BUF U17 ( .A(eCount[14]), .Z(remStepPO[14]));
Q_BUF U18 ( .A(eCount[15]), .Z(remStepPO[15]));
Q_BUF U19 ( .A(eCount[16]), .Z(remStepPO[16]));
Q_BUF U20 ( .A(eCount[17]), .Z(remStepPO[17]));
Q_BUF U21 ( .A(eCount[18]), .Z(remStepPO[18]));
Q_BUF U22 ( .A(eCount[19]), .Z(remStepPO[19]));
Q_BUF U23 ( .A(eCount[20]), .Z(remStepPO[20]));
Q_BUF U24 ( .A(eCount[21]), .Z(remStepPO[21]));
Q_BUF U25 ( .A(eCount[22]), .Z(remStepPO[22]));
Q_BUF U26 ( .A(eCount[23]), .Z(remStepPO[23]));
Q_BUF U27 ( .A(eCount[24]), .Z(remStepPO[24]));
Q_BUF U28 ( .A(eCount[25]), .Z(remStepPO[25]));
Q_BUF U29 ( .A(eCount[26]), .Z(remStepPO[26]));
Q_BUF U30 ( .A(eCount[27]), .Z(remStepPO[27]));
Q_BUF U31 ( .A(eCount[28]), .Z(remStepPO[28]));
Q_BUF U32 ( .A(eCount[29]), .Z(remStepPO[29]));
Q_BUF U33 ( .A(eCount[30]), .Z(remStepPO[30]));
Q_BUF U34 ( .A(eCount[31]), .Z(remStepPO[31]));
Q_BUF U35 ( .A(eCount[32]), .Z(remStepPO[32]));
Q_BUF U36 ( .A(eCount[33]), .Z(remStepPO[33]));
Q_BUF U37 ( .A(eCount[34]), .Z(remStepPO[34]));
Q_BUF U38 ( .A(eCount[35]), .Z(remStepPO[35]));
Q_BUF U39 ( .A(eCount[36]), .Z(remStepPO[36]));
Q_BUF U40 ( .A(eCount[37]), .Z(remStepPO[37]));
Q_BUF U41 ( .A(eCount[38]), .Z(remStepPO[38]));
Q_BUF U42 ( .A(eCount[39]), .Z(remStepPO[39]));
Q_BUF U43 ( .A(eCount[40]), .Z(remStepPO[40]));
Q_BUF U44 ( .A(eCount[41]), .Z(remStepPO[41]));
Q_BUF U45 ( .A(eCount[42]), .Z(remStepPO[42]));
Q_BUF U46 ( .A(eCount[43]), .Z(remStepPO[43]));
Q_BUF U47 ( .A(eCount[44]), .Z(remStepPO[44]));
Q_BUF U48 ( .A(eCount[45]), .Z(remStepPO[45]));
Q_BUF U49 ( .A(eCount[46]), .Z(remStepPO[46]));
Q_BUF U50 ( .A(eCount[47]), .Z(remStepPO[47]));
Q_BUF U51 ( .A(eCount[48]), .Z(remStepPO[48]));
Q_BUF U52 ( .A(eCount[49]), .Z(remStepPO[49]));
Q_BUF U53 ( .A(eCount[50]), .Z(remStepPO[50]));
Q_BUF U54 ( .A(eCount[51]), .Z(remStepPO[51]));
Q_BUF U55 ( .A(eCount[52]), .Z(remStepPO[52]));
Q_BUF U56 ( .A(eCount[53]), .Z(remStepPO[53]));
Q_BUF U57 ( .A(eCount[54]), .Z(remStepPO[54]));
Q_BUF U58 ( .A(eCount[55]), .Z(remStepPO[55]));
Q_BUF U59 ( .A(eCount[56]), .Z(remStepPO[56]));
Q_BUF U60 ( .A(eCount[57]), .Z(remStepPO[57]));
Q_BUF U61 ( .A(eCount[58]), .Z(remStepPO[58]));
Q_BUF U62 ( .A(eCount[59]), .Z(remStepPO[59]));
Q_BUF U63 ( .A(eCount[60]), .Z(remStepPO[60]));
Q_BUF U64 ( .A(eCount[61]), .Z(remStepPO[61]));
Q_BUF U65 ( .A(eCount[62]), .Z(remStepPO[62]));
Q_BUF U66 ( .A(eCount[63]), .Z(remStepPO[63]));
Q_ASSIGN U67 ( .B(stopEmuPI), .A(stopEmuPO));
Q_ASSIGN U68 ( .B(callEmuPI), .A(sendPO));
Q_BUF U69 ( .A(n115), .Z(n1));
Q_AN02 U70 ( .A0(n451), .A1(n518), .Z(n519));
Q_FDP0UA U71 ( .D(dummyW), .QTFCLK( ), .Q(dummyR));
Q_FDP0UA U72 ( .D(memWriteCmd), .QTFCLK( ), .Q(_zzmemWriteCmd));
Q_INV U73 ( .A(callEmu), .Z(n517));
Q_NR02 U74 ( .A0(callEmu), .A1(poBusy), .Z(n516));
Q_INV U75 ( .A(n516), .Z(n518));
Q_XOR2 U76 ( .A0(n518), .A1(evfCount[0]), .Z(n515));
Q_FDP0UA U77 ( .D(n515), .QTFCLK( ), .Q(evfCount[0]));
Q_MX02 U78 ( .S(n516), .A0(n328), .A1(evfCount[1]), .Z(n514));
Q_FDP0UA U79 ( .D(n514), .QTFCLK( ), .Q(evfCount[1]));
Q_MX02 U80 ( .S(n516), .A0(n330), .A1(evfCount[2]), .Z(n513));
Q_FDP0UA U81 ( .D(n513), .QTFCLK( ), .Q(evfCount[2]));
Q_MX02 U82 ( .S(n516), .A0(n332), .A1(evfCount[3]), .Z(n512));
Q_FDP0UA U83 ( .D(n512), .QTFCLK( ), .Q(evfCount[3]));
Q_MX02 U84 ( .S(n516), .A0(n334), .A1(evfCount[4]), .Z(n511));
Q_FDP0UA U85 ( .D(n511), .QTFCLK( ), .Q(evfCount[4]));
Q_MX02 U86 ( .S(n516), .A0(n336), .A1(evfCount[5]), .Z(n510));
Q_FDP0UA U87 ( .D(n510), .QTFCLK( ), .Q(evfCount[5]));
Q_MX02 U88 ( .S(n516), .A0(n338), .A1(evfCount[6]), .Z(n509));
Q_FDP0UA U89 ( .D(n509), .QTFCLK( ), .Q(evfCount[6]));
Q_MX02 U90 ( .S(n516), .A0(n340), .A1(evfCount[7]), .Z(n508));
Q_FDP0UA U91 ( .D(n508), .QTFCLK( ), .Q(evfCount[7]));
Q_MX02 U92 ( .S(n516), .A0(n342), .A1(evfCount[8]), .Z(n507));
Q_FDP0UA U93 ( .D(n507), .QTFCLK( ), .Q(evfCount[8]));
Q_MX02 U94 ( .S(n516), .A0(n344), .A1(evfCount[9]), .Z(n506));
Q_FDP0UA U95 ( .D(n506), .QTFCLK( ), .Q(evfCount[9]));
Q_MX02 U96 ( .S(n516), .A0(n346), .A1(evfCount[10]), .Z(n505));
Q_FDP0UA U97 ( .D(n505), .QTFCLK( ), .Q(evfCount[10]));
Q_MX02 U98 ( .S(n516), .A0(n348), .A1(evfCount[11]), .Z(n504));
Q_FDP0UA U99 ( .D(n504), .QTFCLK( ), .Q(evfCount[11]));
Q_MX02 U100 ( .S(n516), .A0(n350), .A1(evfCount[12]), .Z(n503));
Q_FDP0UA U101 ( .D(n503), .QTFCLK( ), .Q(evfCount[12]));
Q_MX02 U102 ( .S(n516), .A0(n352), .A1(evfCount[13]), .Z(n502));
Q_FDP0UA U103 ( .D(n502), .QTFCLK( ), .Q(evfCount[13]));
Q_MX02 U104 ( .S(n516), .A0(n354), .A1(evfCount[14]), .Z(n501));
Q_FDP0UA U105 ( .D(n501), .QTFCLK( ), .Q(evfCount[14]));
Q_MX02 U106 ( .S(n516), .A0(n356), .A1(evfCount[15]), .Z(n500));
Q_FDP0UA U107 ( .D(n500), .QTFCLK( ), .Q(evfCount[15]));
Q_MX02 U108 ( .S(n516), .A0(n358), .A1(evfCount[16]), .Z(n499));
Q_FDP0UA U109 ( .D(n499), .QTFCLK( ), .Q(evfCount[16]));
Q_MX02 U110 ( .S(n516), .A0(n360), .A1(evfCount[17]), .Z(n498));
Q_FDP0UA U111 ( .D(n498), .QTFCLK( ), .Q(evfCount[17]));
Q_MX02 U112 ( .S(n516), .A0(n362), .A1(evfCount[18]), .Z(n497));
Q_FDP0UA U113 ( .D(n497), .QTFCLK( ), .Q(evfCount[18]));
Q_MX02 U114 ( .S(n516), .A0(n364), .A1(evfCount[19]), .Z(n496));
Q_FDP0UA U115 ( .D(n496), .QTFCLK( ), .Q(evfCount[19]));
Q_MX02 U116 ( .S(n516), .A0(n366), .A1(evfCount[20]), .Z(n495));
Q_FDP0UA U117 ( .D(n495), .QTFCLK( ), .Q(evfCount[20]));
Q_MX02 U118 ( .S(n516), .A0(n368), .A1(evfCount[21]), .Z(n494));
Q_FDP0UA U119 ( .D(n494), .QTFCLK( ), .Q(evfCount[21]));
Q_MX02 U120 ( .S(n516), .A0(n370), .A1(evfCount[22]), .Z(n493));
Q_FDP0UA U121 ( .D(n493), .QTFCLK( ), .Q(evfCount[22]));
Q_MX02 U122 ( .S(n516), .A0(n372), .A1(evfCount[23]), .Z(n492));
Q_FDP0UA U123 ( .D(n492), .QTFCLK( ), .Q(evfCount[23]));
Q_MX02 U124 ( .S(n516), .A0(n374), .A1(evfCount[24]), .Z(n491));
Q_FDP0UA U125 ( .D(n491), .QTFCLK( ), .Q(evfCount[24]));
Q_MX02 U126 ( .S(n516), .A0(n376), .A1(evfCount[25]), .Z(n490));
Q_FDP0UA U127 ( .D(n490), .QTFCLK( ), .Q(evfCount[25]));
Q_MX02 U128 ( .S(n516), .A0(n378), .A1(evfCount[26]), .Z(n489));
Q_FDP0UA U129 ( .D(n489), .QTFCLK( ), .Q(evfCount[26]));
Q_MX02 U130 ( .S(n516), .A0(n380), .A1(evfCount[27]), .Z(n488));
Q_FDP0UA U131 ( .D(n488), .QTFCLK( ), .Q(evfCount[27]));
Q_MX02 U132 ( .S(n516), .A0(n382), .A1(evfCount[28]), .Z(n487));
Q_FDP0UA U133 ( .D(n487), .QTFCLK( ), .Q(evfCount[28]));
Q_MX02 U134 ( .S(n516), .A0(n384), .A1(evfCount[29]), .Z(n486));
Q_FDP0UA U135 ( .D(n486), .QTFCLK( ), .Q(evfCount[29]));
Q_MX02 U136 ( .S(n516), .A0(n386), .A1(evfCount[30]), .Z(n485));
Q_FDP0UA U137 ( .D(n485), .QTFCLK( ), .Q(evfCount[30]));
Q_MX02 U138 ( .S(n516), .A0(n388), .A1(evfCount[31]), .Z(n484));
Q_FDP0UA U139 ( .D(n484), .QTFCLK( ), .Q(evfCount[31]));
Q_MX02 U140 ( .S(n516), .A0(n390), .A1(evfCount[32]), .Z(n483));
Q_FDP0UA U141 ( .D(n483), .QTFCLK( ), .Q(evfCount[32]));
Q_MX02 U142 ( .S(n516), .A0(n392), .A1(evfCount[33]), .Z(n482));
Q_FDP0UA U143 ( .D(n482), .QTFCLK( ), .Q(evfCount[33]));
Q_MX02 U144 ( .S(n516), .A0(n394), .A1(evfCount[34]), .Z(n481));
Q_FDP0UA U145 ( .D(n481), .QTFCLK( ), .Q(evfCount[34]));
Q_MX02 U146 ( .S(n516), .A0(n396), .A1(evfCount[35]), .Z(n480));
Q_FDP0UA U147 ( .D(n480), .QTFCLK( ), .Q(evfCount[35]));
Q_MX02 U148 ( .S(n516), .A0(n398), .A1(evfCount[36]), .Z(n479));
Q_FDP0UA U149 ( .D(n479), .QTFCLK( ), .Q(evfCount[36]));
Q_MX02 U150 ( .S(n516), .A0(n400), .A1(evfCount[37]), .Z(n478));
Q_FDP0UA U151 ( .D(n478), .QTFCLK( ), .Q(evfCount[37]));
Q_MX02 U152 ( .S(n516), .A0(n402), .A1(evfCount[38]), .Z(n477));
Q_FDP0UA U153 ( .D(n477), .QTFCLK( ), .Q(evfCount[38]));
Q_MX02 U154 ( .S(n516), .A0(n404), .A1(evfCount[39]), .Z(n476));
Q_FDP0UA U155 ( .D(n476), .QTFCLK( ), .Q(evfCount[39]));
Q_MX02 U156 ( .S(n516), .A0(n406), .A1(evfCount[40]), .Z(n475));
Q_FDP0UA U157 ( .D(n475), .QTFCLK( ), .Q(evfCount[40]));
Q_MX02 U158 ( .S(n516), .A0(n408), .A1(evfCount[41]), .Z(n474));
Q_FDP0UA U159 ( .D(n474), .QTFCLK( ), .Q(evfCount[41]));
Q_MX02 U160 ( .S(n516), .A0(n410), .A1(evfCount[42]), .Z(n473));
Q_FDP0UA U161 ( .D(n473), .QTFCLK( ), .Q(evfCount[42]));
Q_MX02 U162 ( .S(n516), .A0(n412), .A1(evfCount[43]), .Z(n472));
Q_FDP0UA U163 ( .D(n472), .QTFCLK( ), .Q(evfCount[43]));
Q_MX02 U164 ( .S(n516), .A0(n414), .A1(evfCount[44]), .Z(n471));
Q_FDP0UA U165 ( .D(n471), .QTFCLK( ), .Q(evfCount[44]));
Q_MX02 U166 ( .S(n516), .A0(n416), .A1(evfCount[45]), .Z(n470));
Q_FDP0UA U167 ( .D(n470), .QTFCLK( ), .Q(evfCount[45]));
Q_MX02 U168 ( .S(n516), .A0(n418), .A1(evfCount[46]), .Z(n469));
Q_FDP0UA U169 ( .D(n469), .QTFCLK( ), .Q(evfCount[46]));
Q_MX02 U170 ( .S(n516), .A0(n420), .A1(evfCount[47]), .Z(n468));
Q_FDP0UA U171 ( .D(n468), .QTFCLK( ), .Q(evfCount[47]));
Q_MX02 U172 ( .S(n516), .A0(n422), .A1(evfCount[48]), .Z(n467));
Q_FDP0UA U173 ( .D(n467), .QTFCLK( ), .Q(evfCount[48]));
Q_MX02 U174 ( .S(n516), .A0(n424), .A1(evfCount[49]), .Z(n466));
Q_FDP0UA U175 ( .D(n466), .QTFCLK( ), .Q(evfCount[49]));
Q_MX02 U176 ( .S(n516), .A0(n426), .A1(evfCount[50]), .Z(n465));
Q_FDP0UA U177 ( .D(n465), .QTFCLK( ), .Q(evfCount[50]));
Q_MX02 U178 ( .S(n516), .A0(n428), .A1(evfCount[51]), .Z(n464));
Q_FDP0UA U179 ( .D(n464), .QTFCLK( ), .Q(evfCount[51]));
Q_MX02 U180 ( .S(n516), .A0(n430), .A1(evfCount[52]), .Z(n463));
Q_FDP0UA U181 ( .D(n463), .QTFCLK( ), .Q(evfCount[52]));
Q_MX02 U182 ( .S(n516), .A0(n432), .A1(evfCount[53]), .Z(n462));
Q_FDP0UA U183 ( .D(n462), .QTFCLK( ), .Q(evfCount[53]));
Q_MX02 U184 ( .S(n516), .A0(n434), .A1(evfCount[54]), .Z(n461));
Q_FDP0UA U185 ( .D(n461), .QTFCLK( ), .Q(evfCount[54]));
Q_MX02 U186 ( .S(n516), .A0(n436), .A1(evfCount[55]), .Z(n460));
Q_FDP0UA U187 ( .D(n460), .QTFCLK( ), .Q(evfCount[55]));
Q_MX02 U188 ( .S(n516), .A0(n438), .A1(evfCount[56]), .Z(n459));
Q_FDP0UA U189 ( .D(n459), .QTFCLK( ), .Q(evfCount[56]));
Q_MX02 U190 ( .S(n516), .A0(n440), .A1(evfCount[57]), .Z(n458));
Q_FDP0UA U191 ( .D(n458), .QTFCLK( ), .Q(evfCount[57]));
Q_MX02 U192 ( .S(n516), .A0(n442), .A1(evfCount[58]), .Z(n457));
Q_FDP0UA U193 ( .D(n457), .QTFCLK( ), .Q(evfCount[58]));
Q_MX02 U194 ( .S(n516), .A0(n444), .A1(evfCount[59]), .Z(n456));
Q_FDP0UA U195 ( .D(n456), .QTFCLK( ), .Q(evfCount[59]));
Q_MX02 U196 ( .S(n516), .A0(n446), .A1(evfCount[60]), .Z(n455));
Q_FDP0UA U197 ( .D(n455), .QTFCLK( ), .Q(evfCount[60]));
Q_MX02 U198 ( .S(n516), .A0(n448), .A1(evfCount[61]), .Z(n454));
Q_FDP0UA U199 ( .D(n454), .QTFCLK( ), .Q(evfCount[61]));
Q_MX02 U200 ( .S(n516), .A0(n450), .A1(evfCount[62]), .Z(n453));
Q_FDP0UA U201 ( .D(n453), .QTFCLK( ), .Q(evfCount[62]));
Q_FDP0UA U202 ( .D(n452), .QTFCLK( ), .Q(evfCount[63]));
Q_XOR2 U203 ( .A0(evfCount[63]), .A1(n519), .Z(n452));
Q_AD01HF U204 ( .A0(evfCount[62]), .B0(n449), .S(n450), .CO(n451));
Q_AD01HF U205 ( .A0(evfCount[61]), .B0(n447), .S(n448), .CO(n449));
Q_AD01HF U206 ( .A0(evfCount[60]), .B0(n445), .S(n446), .CO(n447));
Q_AD01HF U207 ( .A0(evfCount[59]), .B0(n443), .S(n444), .CO(n445));
Q_AD01HF U208 ( .A0(evfCount[58]), .B0(n441), .S(n442), .CO(n443));
Q_AD01HF U209 ( .A0(evfCount[57]), .B0(n439), .S(n440), .CO(n441));
Q_AD01HF U210 ( .A0(evfCount[56]), .B0(n437), .S(n438), .CO(n439));
Q_AD01HF U211 ( .A0(evfCount[55]), .B0(n435), .S(n436), .CO(n437));
Q_AD01HF U212 ( .A0(evfCount[54]), .B0(n433), .S(n434), .CO(n435));
Q_AD01HF U213 ( .A0(evfCount[53]), .B0(n431), .S(n432), .CO(n433));
Q_AD01HF U214 ( .A0(evfCount[52]), .B0(n429), .S(n430), .CO(n431));
Q_AD01HF U215 ( .A0(evfCount[51]), .B0(n427), .S(n428), .CO(n429));
Q_AD01HF U216 ( .A0(evfCount[50]), .B0(n425), .S(n426), .CO(n427));
Q_AD01HF U217 ( .A0(evfCount[49]), .B0(n423), .S(n424), .CO(n425));
Q_AD01HF U218 ( .A0(evfCount[48]), .B0(n421), .S(n422), .CO(n423));
Q_AD01HF U219 ( .A0(evfCount[47]), .B0(n419), .S(n420), .CO(n421));
Q_AD01HF U220 ( .A0(evfCount[46]), .B0(n417), .S(n418), .CO(n419));
Q_AD01HF U221 ( .A0(evfCount[45]), .B0(n415), .S(n416), .CO(n417));
Q_AD01HF U222 ( .A0(evfCount[44]), .B0(n413), .S(n414), .CO(n415));
Q_AD01HF U223 ( .A0(evfCount[43]), .B0(n411), .S(n412), .CO(n413));
Q_AD01HF U224 ( .A0(evfCount[42]), .B0(n409), .S(n410), .CO(n411));
Q_AD01HF U225 ( .A0(evfCount[41]), .B0(n407), .S(n408), .CO(n409));
Q_AD01HF U226 ( .A0(evfCount[40]), .B0(n405), .S(n406), .CO(n407));
Q_AD01HF U227 ( .A0(evfCount[39]), .B0(n403), .S(n404), .CO(n405));
Q_AD01HF U228 ( .A0(evfCount[38]), .B0(n401), .S(n402), .CO(n403));
Q_AD01HF U229 ( .A0(evfCount[37]), .B0(n399), .S(n400), .CO(n401));
Q_AD01HF U230 ( .A0(evfCount[36]), .B0(n397), .S(n398), .CO(n399));
Q_AD01HF U231 ( .A0(evfCount[35]), .B0(n395), .S(n396), .CO(n397));
Q_AD01HF U232 ( .A0(evfCount[34]), .B0(n393), .S(n394), .CO(n395));
Q_AD01HF U233 ( .A0(evfCount[33]), .B0(n391), .S(n392), .CO(n393));
Q_AD01HF U234 ( .A0(evfCount[32]), .B0(n389), .S(n390), .CO(n391));
Q_AD01HF U235 ( .A0(evfCount[31]), .B0(n387), .S(n388), .CO(n389));
Q_AD01HF U236 ( .A0(evfCount[30]), .B0(n385), .S(n386), .CO(n387));
Q_AD01HF U237 ( .A0(evfCount[29]), .B0(n383), .S(n384), .CO(n385));
Q_AD01HF U238 ( .A0(evfCount[28]), .B0(n381), .S(n382), .CO(n383));
Q_AD01HF U239 ( .A0(evfCount[27]), .B0(n379), .S(n380), .CO(n381));
Q_AD01HF U240 ( .A0(evfCount[26]), .B0(n377), .S(n378), .CO(n379));
Q_AD01HF U241 ( .A0(evfCount[25]), .B0(n375), .S(n376), .CO(n377));
Q_AD01HF U242 ( .A0(evfCount[24]), .B0(n373), .S(n374), .CO(n375));
Q_AD01HF U243 ( .A0(evfCount[23]), .B0(n371), .S(n372), .CO(n373));
Q_AD01HF U244 ( .A0(evfCount[22]), .B0(n369), .S(n370), .CO(n371));
Q_AD01HF U245 ( .A0(evfCount[21]), .B0(n367), .S(n368), .CO(n369));
Q_AD01HF U246 ( .A0(evfCount[20]), .B0(n365), .S(n366), .CO(n367));
Q_AD01HF U247 ( .A0(evfCount[19]), .B0(n363), .S(n364), .CO(n365));
Q_AD01HF U248 ( .A0(evfCount[18]), .B0(n361), .S(n362), .CO(n363));
Q_AD01HF U249 ( .A0(evfCount[17]), .B0(n359), .S(n360), .CO(n361));
Q_AD01HF U250 ( .A0(evfCount[16]), .B0(n357), .S(n358), .CO(n359));
Q_AD01HF U251 ( .A0(evfCount[15]), .B0(n355), .S(n356), .CO(n357));
Q_AD01HF U252 ( .A0(evfCount[14]), .B0(n353), .S(n354), .CO(n355));
Q_AD01HF U253 ( .A0(evfCount[13]), .B0(n351), .S(n352), .CO(n353));
Q_AD01HF U254 ( .A0(evfCount[12]), .B0(n349), .S(n350), .CO(n351));
Q_AD01HF U255 ( .A0(evfCount[11]), .B0(n347), .S(n348), .CO(n349));
Q_AD01HF U256 ( .A0(evfCount[10]), .B0(n345), .S(n346), .CO(n347));
Q_AD01HF U257 ( .A0(evfCount[9]), .B0(n343), .S(n344), .CO(n345));
Q_AD01HF U258 ( .A0(evfCount[8]), .B0(n341), .S(n342), .CO(n343));
Q_AD01HF U259 ( .A0(evfCount[7]), .B0(n339), .S(n340), .CO(n341));
Q_AD01HF U260 ( .A0(evfCount[6]), .B0(n337), .S(n338), .CO(n339));
Q_AD01HF U261 ( .A0(evfCount[5]), .B0(n335), .S(n336), .CO(n337));
Q_AD01HF U262 ( .A0(evfCount[4]), .B0(n333), .S(n334), .CO(n335));
Q_AD01HF U263 ( .A0(evfCount[3]), .B0(n331), .S(n332), .CO(n333));
Q_AD01HF U264 ( .A0(evfCount[2]), .B0(n329), .S(n330), .CO(n331));
Q_AD01HF U265 ( .A0(evfCount[1]), .B0(evfCount[0]), .S(n328), .CO(n329));
Q_NR02 U266 ( .A0(callEmu), .A1(n327), .Z(n326));
Q_MX02 U267 ( .S(n326), .A0(n310), .A1(evalOnDExt[0]), .Z(n325));
Q_FDP0UA U268 ( .D(n325), .QTFCLK( ), .Q(evalOnDExt[0]));
Q_MX02 U269 ( .S(n326), .A0(n311), .A1(evalOnDExt[1]), .Z(n324));
Q_FDP0UA U270 ( .D(n324), .QTFCLK( ), .Q(evalOnDExt[1]));
Q_MX02 U271 ( .S(n326), .A0(n312), .A1(evalOnDExt[2]), .Z(n323));
Q_FDP0UA U272 ( .D(n323), .QTFCLK( ), .Q(evalOnDExt[2]));
Q_MX02 U273 ( .S(n326), .A0(n313), .A1(evalOnDExt[3]), .Z(n322));
Q_FDP0UA U274 ( .D(n322), .QTFCLK( ), .Q(evalOnDExt[3]));
Q_MX02 U275 ( .S(n326), .A0(n314), .A1(evalOnDExt[4]), .Z(n321));
Q_FDP0UA U276 ( .D(n321), .QTFCLK( ), .Q(evalOnDExt[4]));
Q_MX02 U277 ( .S(n326), .A0(n315), .A1(evalOnDExt[5]), .Z(n320));
Q_FDP0UA U278 ( .D(n320), .QTFCLK( ), .Q(evalOnDExt[5]));
Q_MX02 U279 ( .S(n326), .A0(n316), .A1(evalOnDExt[6]), .Z(n319));
Q_FDP0UA U280 ( .D(n319), .QTFCLK( ), .Q(evalOnDExt[6]));
Q_MX02 U281 ( .S(n326), .A0(n317), .A1(evalOnDExt[7]), .Z(n318));
Q_FDP0UA U282 ( .D(n318), .QTFCLK( ), .Q(evalOnDExt[7]));
Q_FDP0UA U283 ( .D(n292), .QTFCLK( ), .Q(callEmuD));
Q_MX02 U284 ( .S(callEmu), .A0(n309), .A1(evalOnDCtl[7]), .Z(n317));
Q_MX02 U285 ( .S(callEmu), .A0(n307), .A1(evalOnDCtl[6]), .Z(n316));
Q_MX02 U286 ( .S(callEmu), .A0(n305), .A1(evalOnDCtl[5]), .Z(n315));
Q_MX02 U287 ( .S(callEmu), .A0(n303), .A1(evalOnDCtl[4]), .Z(n314));
Q_MX02 U288 ( .S(callEmu), .A0(n301), .A1(evalOnDCtl[3]), .Z(n313));
Q_MX02 U289 ( .S(callEmu), .A0(n299), .A1(evalOnDCtl[2]), .Z(n312));
Q_MX02 U290 ( .S(callEmu), .A0(n297), .A1(evalOnDCtl[1]), .Z(n311));
Q_MX02 U291 ( .S(callEmu), .A0(n296), .A1(evalOnDCtl[0]), .Z(n310));
Q_XNR2 U292 ( .A0(evalOnDExt[7]), .A1(n308), .Z(n309));
Q_OR02 U293 ( .A0(evalOnDExt[6]), .A1(n306), .Z(n308));
Q_XNR2 U294 ( .A0(evalOnDExt[6]), .A1(n306), .Z(n307));
Q_OR02 U295 ( .A0(evalOnDExt[5]), .A1(n304), .Z(n306));
Q_XNR2 U296 ( .A0(evalOnDExt[5]), .A1(n304), .Z(n305));
Q_OR02 U297 ( .A0(evalOnDExt[4]), .A1(n302), .Z(n304));
Q_XNR2 U298 ( .A0(evalOnDExt[4]), .A1(n302), .Z(n303));
Q_OR02 U299 ( .A0(evalOnDExt[3]), .A1(n300), .Z(n302));
Q_XNR2 U300 ( .A0(evalOnDExt[3]), .A1(n300), .Z(n301));
Q_OR02 U301 ( .A0(evalOnDExt[2]), .A1(n298), .Z(n300));
Q_XNR2 U302 ( .A0(evalOnDExt[2]), .A1(n298), .Z(n299));
Q_OR02 U303 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .Z(n298));
Q_XNR2 U304 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .Z(n297));
Q_INV U305 ( .A(evalOnDExt[0]), .Z(n296));
Q_OR02 U306 ( .A0(n294), .A1(n295), .Z(n327));
Q_OR03 U307 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .A2(n293), .Z(n295));
Q_OR03 U308 ( .A0(evalOnDExt[4]), .A1(evalOnDExt[3]), .A2(evalOnDExt[2]), .Z(n294));
Q_OR03 U309 ( .A0(evalOnDExt[7]), .A1(evalOnDExt[6]), .A2(evalOnDExt[5]), .Z(n293));
Q_OR02 U310 ( .A0(callEmu), .A1(poBusy), .Z(n292));
Q_FDP0UA U311 ( .D(FvUseOnly), .QTFCLK( ), .Q(FvUseOnlyR));
Q_FDP0UA U312 ( .D(APPLY_PI), .QTFCLK( ), .Q(applyPiR));
Q_FDP0UA U313 ( .D(n284), .QTFCLK( ), .Q(poDelay[0]));
Q_FDP0UA U314 ( .D(n285), .QTFCLK( ), .Q(poDelay[1]));
Q_FDP0UA U315 ( .D(n286), .QTFCLK( ), .Q(poDelay[2]));
Q_FDP0UA U316 ( .D(n287), .QTFCLK( ), .Q(poDelay[3]));
Q_FDP0UA U317 ( .D(n288), .QTFCLK( ), .Q(poDelay[4]));
Q_FDP0UA U318 ( .D(n289), .QTFCLK( ), .Q(poDelay[5]));
Q_FDP0UA U319 ( .D(n290), .QTFCLK( ), .Q(poDelay[6]));
Q_FDP0UA U320 ( .D(n291), .QTFCLK( ), .Q(poDelay[7]));
Q_MX02 U321 ( .S(callEmu), .A0(n283), .A1(fclkPerEval[7]), .Z(n291));
Q_MX02 U322 ( .S(callEmu), .A0(n282), .A1(fclkPerEval[6]), .Z(n290));
Q_MX02 U323 ( .S(callEmu), .A0(n281), .A1(fclkPerEval[5]), .Z(n289));
Q_MX02 U324 ( .S(callEmu), .A0(n280), .A1(fclkPerEval[4]), .Z(n288));
Q_MX02 U325 ( .S(callEmu), .A0(n279), .A1(fclkPerEval[3]), .Z(n287));
Q_MX02 U326 ( .S(callEmu), .A0(n278), .A1(fclkPerEval[2]), .Z(n286));
Q_MX02 U327 ( .S(callEmu), .A0(n277), .A1(fclkPerEval[1]), .Z(n285));
Q_MX02 U328 ( .S(callEmu), .A0(n276), .A1(fclkPerEval[0]), .Z(n284));
Q_AN02 U329 ( .A0(poBusy), .A1(n275), .Z(n283));
Q_AN02 U330 ( .A0(poBusy), .A1(n273), .Z(n282));
Q_AN02 U331 ( .A0(poBusy), .A1(n271), .Z(n281));
Q_AN02 U332 ( .A0(poBusy), .A1(n269), .Z(n280));
Q_AN02 U333 ( .A0(poBusy), .A1(n267), .Z(n279));
Q_AN02 U334 ( .A0(poBusy), .A1(n265), .Z(n278));
Q_AN02 U335 ( .A0(poBusy), .A1(n263), .Z(n277));
Q_AN02 U336 ( .A0(poBusy), .A1(n262), .Z(n276));
Q_XNR2 U337 ( .A0(poDelay[7]), .A1(n274), .Z(n275));
Q_OR02 U338 ( .A0(poDelay[6]), .A1(n272), .Z(n274));
Q_XNR2 U339 ( .A0(poDelay[6]), .A1(n272), .Z(n273));
Q_OR02 U340 ( .A0(poDelay[5]), .A1(n270), .Z(n272));
Q_XNR2 U341 ( .A0(poDelay[5]), .A1(n270), .Z(n271));
Q_OR02 U342 ( .A0(poDelay[4]), .A1(n268), .Z(n270));
Q_XNR2 U343 ( .A0(poDelay[4]), .A1(n268), .Z(n269));
Q_OR02 U344 ( .A0(poDelay[3]), .A1(n266), .Z(n268));
Q_XNR2 U345 ( .A0(poDelay[3]), .A1(n266), .Z(n267));
Q_OR02 U346 ( .A0(poDelay[2]), .A1(n264), .Z(n266));
Q_XNR2 U347 ( .A0(poDelay[2]), .A1(n264), .Z(n265));
Q_OR02 U348 ( .A0(poDelay[1]), .A1(poDelay[0]), .Z(n264));
Q_XNR2 U349 ( .A0(poDelay[1]), .A1(poDelay[0]), .Z(n263));
Q_INV U350 ( .A(poDelay[0]), .Z(n262));
Q_FDP0UA U351 ( .D(lbrOn), .QTFCLK( ), .Q(lbrOnD));
Q_FDP0UA U352 ( .D(sendPO), .QTFCLK( ), .Q(callEmuR));
Q_FDP0UA U353 ( .D(fclkPerEval[7]), .QTFCLK( ), .Q(fclkPerEval[7]));
Q_FDP0UA U354 ( .D(fclkPerEval[6]), .QTFCLK( ), .Q(fclkPerEval[6]));
Q_FDP0UA U355 ( .D(fclkPerEval[5]), .QTFCLK( ), .Q(fclkPerEval[5]));
Q_FDP0UA U356 ( .D(fclkPerEval[4]), .QTFCLK( ), .Q(fclkPerEval[4]));
Q_FDP0UA U357 ( .D(fclkPerEval[3]), .QTFCLK( ), .Q(fclkPerEval[3]));
Q_FDP0UA U358 ( .D(fclkPerEval[2]), .QTFCLK( ), .Q(fclkPerEval[2]));
Q_FDP0UA U359 ( .D(fclkPerEval[1]), .QTFCLK( ), .Q(fclkPerEval[1]));
Q_FDP0UA U360 ( .D(fclkPerEval[0]), .QTFCLK( ), .Q(fclkPerEval[0]));
Q_FDP0UA U361 ( .D(sdlEnable), .QTFCLK( ), .Q(sdlEnable));
Q_FDP0UA U362 ( .D(tbcEnable), .QTFCLK( ), .Q(tbcEnable));
Q_FDP0UA U363 ( .D(evalOnDCtl[7]), .QTFCLK( ), .Q(evalOnDCtl[7]));
Q_FDP0UA U364 ( .D(evalOnDCtl[6]), .QTFCLK( ), .Q(evalOnDCtl[6]));
Q_FDP0UA U365 ( .D(evalOnDCtl[5]), .QTFCLK( ), .Q(evalOnDCtl[5]));
Q_FDP0UA U366 ( .D(evalOnDCtl[4]), .QTFCLK( ), .Q(evalOnDCtl[4]));
Q_FDP0UA U367 ( .D(evalOnDCtl[3]), .QTFCLK( ), .Q(evalOnDCtl[3]));
Q_FDP0UA U368 ( .D(evalOnDCtl[2]), .QTFCLK( ), .Q(evalOnDCtl[2]));
Q_FDP0UA U369 ( .D(evalOnDCtl[1]), .QTFCLK( ), .Q(evalOnDCtl[1]));
Q_FDP0UA U370 ( .D(evalOnDCtl[0]), .QTFCLK( ), .Q(evalOnDCtl[0]));
Q_FDP0UA U371 ( .D(hotSwapOnPI), .QTFCLK( ), .Q(hotSwapOnPI));
Q_FDP0UA U372 ( .D(sdlHaltHwClk), .QTFCLK( ), .Q(sdlHaltHwClk));
Q_FDP0UA U373 ( .D(hwClkDbg), .QTFCLK( ), .Q(hwClkDbg));
Q_FDP0UA U374 ( .D(hwClkDbgTime), .QTFCLK( ), .Q(hwClkDbgTime));
Q_FDP0UA U375 ( .D(hwClkEnable), .QTFCLK( ), .Q(hwClkEnable));
Q_FDP0UA U376 ( .D(gfifoOff), .QTFCLK( ), .Q(gfifoOff));
Q_FDP0UA U377 ( .D(hssReset), .QTFCLK( ), .Q(hssReset));
Q_XOR2 U378 ( .A0(_zzmemWriteCmd), .A1(memWriteCmd), .Z(n260));
Q_BUFZP U379 ( .OE(n260), .A(n259), .Z(asyncCall));
Q_FDP0 eClkR_REG  ( .CK(rClk), .D(eClkv), .Q(eClkR), .QN( ));
Q_AD01HF U381 ( .A0(remStepPO[1]), .B0(remStepPO[0]), .S(n257), .CO(n256));
Q_AD01HF U382 ( .A0(remStepPO[2]), .B0(n256), .S(n255), .CO(n254));
Q_AD01HF U383 ( .A0(remStepPO[3]), .B0(n254), .S(n253), .CO(n252));
Q_AD01HF U384 ( .A0(remStepPO[4]), .B0(n252), .S(n251), .CO(n250));
Q_AD01HF U385 ( .A0(remStepPO[5]), .B0(n250), .S(n249), .CO(n248));
Q_AD01HF U386 ( .A0(remStepPO[6]), .B0(n248), .S(n247), .CO(n246));
Q_AD01HF U387 ( .A0(remStepPO[7]), .B0(n246), .S(n245), .CO(n244));
Q_AD01HF U388 ( .A0(remStepPO[8]), .B0(n244), .S(n243), .CO(n242));
Q_AD01HF U389 ( .A0(remStepPO[9]), .B0(n242), .S(n241), .CO(n240));
Q_AD01HF U390 ( .A0(remStepPO[10]), .B0(n240), .S(n239), .CO(n238));
Q_AD01HF U391 ( .A0(remStepPO[11]), .B0(n238), .S(n237), .CO(n236));
Q_AD01HF U392 ( .A0(remStepPO[12]), .B0(n236), .S(n235), .CO(n234));
Q_AD01HF U393 ( .A0(remStepPO[13]), .B0(n234), .S(n233), .CO(n232));
Q_AD01HF U394 ( .A0(remStepPO[14]), .B0(n232), .S(n231), .CO(n230));
Q_AD01HF U395 ( .A0(remStepPO[15]), .B0(n230), .S(n229), .CO(n228));
Q_AD01HF U396 ( .A0(remStepPO[16]), .B0(n228), .S(n227), .CO(n226));
Q_AD01HF U397 ( .A0(remStepPO[17]), .B0(n226), .S(n225), .CO(n224));
Q_AD01HF U398 ( .A0(remStepPO[18]), .B0(n224), .S(n223), .CO(n222));
Q_AD01HF U399 ( .A0(remStepPO[19]), .B0(n222), .S(n221), .CO(n220));
Q_AD01HF U400 ( .A0(remStepPO[20]), .B0(n220), .S(n219), .CO(n218));
Q_AD01HF U401 ( .A0(remStepPO[21]), .B0(n218), .S(n217), .CO(n216));
Q_AD01HF U402 ( .A0(remStepPO[22]), .B0(n216), .S(n215), .CO(n214));
Q_AD01HF U403 ( .A0(remStepPO[23]), .B0(n214), .S(n213), .CO(n212));
Q_AD01HF U404 ( .A0(remStepPO[24]), .B0(n212), .S(n211), .CO(n210));
Q_AD01HF U405 ( .A0(remStepPO[25]), .B0(n210), .S(n209), .CO(n208));
Q_AD01HF U406 ( .A0(remStepPO[26]), .B0(n208), .S(n207), .CO(n206));
Q_AD01HF U407 ( .A0(remStepPO[27]), .B0(n206), .S(n205), .CO(n204));
Q_AD01HF U408 ( .A0(remStepPO[28]), .B0(n204), .S(n203), .CO(n202));
Q_AD01HF U409 ( .A0(remStepPO[29]), .B0(n202), .S(n201), .CO(n200));
Q_AD01HF U410 ( .A0(remStepPO[30]), .B0(n200), .S(n199), .CO(n198));
Q_AD01HF U411 ( .A0(remStepPO[31]), .B0(n198), .S(n197), .CO(n196));
Q_AD01HF U412 ( .A0(remStepPO[32]), .B0(n196), .S(n195), .CO(n194));
Q_AD01HF U413 ( .A0(remStepPO[33]), .B0(n194), .S(n193), .CO(n192));
Q_AD01HF U414 ( .A0(remStepPO[34]), .B0(n192), .S(n191), .CO(n190));
Q_AD01HF U415 ( .A0(remStepPO[35]), .B0(n190), .S(n189), .CO(n188));
Q_AD01HF U416 ( .A0(remStepPO[36]), .B0(n188), .S(n187), .CO(n186));
Q_AD01HF U417 ( .A0(remStepPO[37]), .B0(n186), .S(n185), .CO(n184));
Q_AD01HF U418 ( .A0(remStepPO[38]), .B0(n184), .S(n183), .CO(n182));
Q_AD01HF U419 ( .A0(remStepPO[39]), .B0(n182), .S(n181), .CO(n180));
Q_AD01HF U420 ( .A0(remStepPO[40]), .B0(n180), .S(n179), .CO(n178));
Q_AD01HF U421 ( .A0(remStepPO[41]), .B0(n178), .S(n177), .CO(n176));
Q_AD01HF U422 ( .A0(remStepPO[42]), .B0(n176), .S(n175), .CO(n174));
Q_AD01HF U423 ( .A0(remStepPO[43]), .B0(n174), .S(n173), .CO(n172));
Q_AD01HF U424 ( .A0(remStepPO[44]), .B0(n172), .S(n171), .CO(n170));
Q_AD01HF U425 ( .A0(remStepPO[45]), .B0(n170), .S(n169), .CO(n168));
Q_AD01HF U426 ( .A0(remStepPO[46]), .B0(n168), .S(n167), .CO(n166));
Q_AD01HF U427 ( .A0(remStepPO[47]), .B0(n166), .S(n165), .CO(n164));
Q_AD01HF U428 ( .A0(remStepPO[48]), .B0(n164), .S(n163), .CO(n162));
Q_AD01HF U429 ( .A0(remStepPO[49]), .B0(n162), .S(n161), .CO(n160));
Q_AD01HF U430 ( .A0(remStepPO[50]), .B0(n160), .S(n159), .CO(n158));
Q_AD01HF U431 ( .A0(remStepPO[51]), .B0(n158), .S(n157), .CO(n156));
Q_AD01HF U432 ( .A0(remStepPO[52]), .B0(n156), .S(n155), .CO(n154));
Q_AD01HF U433 ( .A0(remStepPO[53]), .B0(n154), .S(n153), .CO(n152));
Q_AD01HF U434 ( .A0(remStepPO[54]), .B0(n152), .S(n151), .CO(n150));
Q_AD01HF U435 ( .A0(remStepPO[55]), .B0(n150), .S(n149), .CO(n148));
Q_AD01HF U436 ( .A0(remStepPO[56]), .B0(n148), .S(n147), .CO(n146));
Q_AD01HF U437 ( .A0(remStepPO[57]), .B0(n146), .S(n145), .CO(n144));
Q_AD01HF U438 ( .A0(remStepPO[58]), .B0(n144), .S(n143), .CO(n142));
Q_AD01HF U439 ( .A0(remStepPO[59]), .B0(n142), .S(n141), .CO(n140));
Q_AD01HF U440 ( .A0(remStepPO[60]), .B0(n140), .S(n139), .CO(n138));
Q_AD01HF U441 ( .A0(remStepPO[61]), .B0(n138), .S(n137), .CO(n136));
Q_AD01HF U442 ( .A0(remStepPO[62]), .B0(n136), .S(n135), .CO(n134));
Q_FDP0 \eCount_REG[62] ( .CK(rClk), .D(n135), .Q(eCount[62]), .QN( ));
Q_FDP0 \eCount_REG[61] ( .CK(rClk), .D(n137), .Q(eCount[61]), .QN( ));
Q_FDP0 \eCount_REG[60] ( .CK(rClk), .D(n139), .Q(eCount[60]), .QN( ));
Q_FDP0 \eCount_REG[59] ( .CK(rClk), .D(n141), .Q(eCount[59]), .QN( ));
Q_FDP0 \eCount_REG[58] ( .CK(rClk), .D(n143), .Q(eCount[58]), .QN( ));
Q_FDP0 \eCount_REG[57] ( .CK(rClk), .D(n145), .Q(eCount[57]), .QN( ));
Q_FDP0 \eCount_REG[56] ( .CK(rClk), .D(n147), .Q(eCount[56]), .QN( ));
Q_FDP0 \eCount_REG[55] ( .CK(rClk), .D(n149), .Q(eCount[55]), .QN( ));
Q_FDP0 \eCount_REG[54] ( .CK(rClk), .D(n151), .Q(eCount[54]), .QN( ));
Q_FDP0 \eCount_REG[53] ( .CK(rClk), .D(n153), .Q(eCount[53]), .QN( ));
Q_FDP0 \eCount_REG[52] ( .CK(rClk), .D(n155), .Q(eCount[52]), .QN( ));
Q_FDP0 \eCount_REG[51] ( .CK(rClk), .D(n157), .Q(eCount[51]), .QN( ));
Q_FDP0 \eCount_REG[50] ( .CK(rClk), .D(n159), .Q(eCount[50]), .QN( ));
Q_FDP0 \eCount_REG[49] ( .CK(rClk), .D(n161), .Q(eCount[49]), .QN( ));
Q_FDP0 \eCount_REG[48] ( .CK(rClk), .D(n163), .Q(eCount[48]), .QN( ));
Q_FDP0 \eCount_REG[47] ( .CK(rClk), .D(n165), .Q(eCount[47]), .QN( ));
Q_FDP0 \eCount_REG[46] ( .CK(rClk), .D(n167), .Q(eCount[46]), .QN( ));
Q_FDP0 \eCount_REG[45] ( .CK(rClk), .D(n169), .Q(eCount[45]), .QN( ));
Q_FDP0 \eCount_REG[44] ( .CK(rClk), .D(n171), .Q(eCount[44]), .QN( ));
Q_FDP0 \eCount_REG[43] ( .CK(rClk), .D(n173), .Q(eCount[43]), .QN( ));
Q_FDP0 \eCount_REG[42] ( .CK(rClk), .D(n175), .Q(eCount[42]), .QN( ));
Q_FDP0 \eCount_REG[41] ( .CK(rClk), .D(n177), .Q(eCount[41]), .QN( ));
Q_FDP0 \eCount_REG[40] ( .CK(rClk), .D(n179), .Q(eCount[40]), .QN( ));
Q_FDP0 \eCount_REG[39] ( .CK(rClk), .D(n181), .Q(eCount[39]), .QN( ));
Q_FDP0 \eCount_REG[38] ( .CK(rClk), .D(n183), .Q(eCount[38]), .QN( ));
Q_FDP0 \eCount_REG[37] ( .CK(rClk), .D(n185), .Q(eCount[37]), .QN( ));
Q_FDP0 \eCount_REG[36] ( .CK(rClk), .D(n187), .Q(eCount[36]), .QN( ));
Q_FDP0 \eCount_REG[35] ( .CK(rClk), .D(n189), .Q(eCount[35]), .QN( ));
Q_FDP0 \eCount_REG[34] ( .CK(rClk), .D(n191), .Q(eCount[34]), .QN( ));
Q_FDP0 \eCount_REG[33] ( .CK(rClk), .D(n193), .Q(eCount[33]), .QN( ));
Q_FDP0 \eCount_REG[32] ( .CK(rClk), .D(n195), .Q(eCount[32]), .QN( ));
Q_FDP0 \eCount_REG[31] ( .CK(rClk), .D(n197), .Q(eCount[31]), .QN( ));
Q_FDP0 \eCount_REG[30] ( .CK(rClk), .D(n199), .Q(eCount[30]), .QN( ));
Q_FDP0 \eCount_REG[29] ( .CK(rClk), .D(n201), .Q(eCount[29]), .QN( ));
Q_FDP0 \eCount_REG[28] ( .CK(rClk), .D(n203), .Q(eCount[28]), .QN( ));
Q_FDP0 \eCount_REG[27] ( .CK(rClk), .D(n205), .Q(eCount[27]), .QN( ));
Q_FDP0 \eCount_REG[26] ( .CK(rClk), .D(n207), .Q(eCount[26]), .QN( ));
Q_FDP0 \eCount_REG[25] ( .CK(rClk), .D(n209), .Q(eCount[25]), .QN( ));
Q_FDP0 \eCount_REG[24] ( .CK(rClk), .D(n211), .Q(eCount[24]), .QN( ));
Q_FDP0 \eCount_REG[23] ( .CK(rClk), .D(n213), .Q(eCount[23]), .QN( ));
Q_FDP0 \eCount_REG[22] ( .CK(rClk), .D(n215), .Q(eCount[22]), .QN( ));
Q_FDP0 \eCount_REG[21] ( .CK(rClk), .D(n217), .Q(eCount[21]), .QN( ));
Q_FDP0 \eCount_REG[20] ( .CK(rClk), .D(n219), .Q(eCount[20]), .QN( ));
Q_FDP0 \eCount_REG[19] ( .CK(rClk), .D(n221), .Q(eCount[19]), .QN( ));
Q_FDP0 \eCount_REG[18] ( .CK(rClk), .D(n223), .Q(eCount[18]), .QN( ));
Q_FDP0 \eCount_REG[17] ( .CK(rClk), .D(n225), .Q(eCount[17]), .QN( ));
Q_FDP0 \eCount_REG[16] ( .CK(rClk), .D(n227), .Q(eCount[16]), .QN( ));
Q_FDP0 \eCount_REG[15] ( .CK(rClk), .D(n229), .Q(eCount[15]), .QN( ));
Q_FDP0 \eCount_REG[14] ( .CK(rClk), .D(n231), .Q(eCount[14]), .QN( ));
Q_FDP0 \eCount_REG[13] ( .CK(rClk), .D(n233), .Q(eCount[13]), .QN( ));
Q_FDP0 \eCount_REG[12] ( .CK(rClk), .D(n235), .Q(eCount[12]), .QN( ));
Q_FDP0 \eCount_REG[11] ( .CK(rClk), .D(n237), .Q(eCount[11]), .QN( ));
Q_FDP0 \eCount_REG[10] ( .CK(rClk), .D(n239), .Q(eCount[10]), .QN( ));
Q_FDP0 \eCount_REG[9] ( .CK(rClk), .D(n241), .Q(eCount[9]), .QN( ));
Q_FDP0 \eCount_REG[8] ( .CK(rClk), .D(n243), .Q(eCount[8]), .QN( ));
Q_FDP0 \eCount_REG[7] ( .CK(rClk), .D(n245), .Q(eCount[7]), .QN( ));
Q_FDP0 \eCount_REG[6] ( .CK(rClk), .D(n247), .Q(eCount[6]), .QN( ));
Q_FDP0 \eCount_REG[5] ( .CK(rClk), .D(n249), .Q(eCount[5]), .QN( ));
Q_FDP0 \eCount_REG[4] ( .CK(rClk), .D(n251), .Q(eCount[4]), .QN( ));
Q_FDP0 \eCount_REG[3] ( .CK(rClk), .D(n253), .Q(eCount[3]), .QN( ));
Q_FDP0 \eCount_REG[2] ( .CK(rClk), .D(n255), .Q(eCount[2]), .QN( ));
Q_FDP0 \eCount_REG[1] ( .CK(rClk), .D(n257), .Q(eCount[1]), .QN( ));
Q_FDP0 \eCount_REG[0] ( .CK(rClk), .D(n258), .Q(eCount[0]), .QN(n258));
Q_LDP0 stopCPFPO_REG  ( .G(callEmu), .D(cpfStop), .Q(stopCPFPO), .QN( ));
Q_LDP0 stopSDLPO_REG  ( .G(callEmu), .D(n127), .Q(stopSDLPO), .QN( ));
Q_AN02 U508 ( .A0(dbiEvent), .A1(n517), .Z(FvUseOnly));
Q_OR02 U509 ( .A0(lbrOn), .A1(lbrOnD), .Z(evalOn));
Q_LDP0 stop3PO_REG  ( .G(callEmu), .D(n133), .Q(stop3PO), .QN( ));
Q_OR03 U511 ( .A0(stopEmuPO), .A1(n127), .A2(cpfStop), .Z(n133));
Q_LDP0 stop4PO_REG  ( .G(callEmu), .D(n126), .Q(stop4PO), .QN( ));
Q_LDP0 stop2PO_REG  ( .G(callEmu), .D(n125), .Q(stop2PO), .QN( ));
Q_LDP0 stop1PO_REG  ( .G(callEmu), .D(n124), .Q(stop1PO), .QN( ));
Q_NR03 U515 ( .A0(n132), .A1(poDelay[1]), .A2(n131), .Z(tbcPO));
Q_OR02 U516 ( .A0(poDelay[3]), .A1(poDelay[2]), .Z(n132));
Q_OR03 U517 ( .A0(poDelay[7]), .A1(poDelay[6]), .A2(n130), .Z(n131));
Q_OR02 U518 ( .A0(poDelay[5]), .A1(poDelay[4]), .Z(n130));
Q_OR03 U519 ( .A0(evalOnOrig), .A1(n327), .A2(asyncCall), .Z(lbrOn));
Q_OR02 U520 ( .A0(callEmu), .A1(hotSwapOnPI), .Z(eventOn));
Q_OR02 U521 ( .A0(callEmu), .A1(n129), .Z(evalOnOrig));
Q_OR03 U522 ( .A0(bWait), .A1(callEmuD), .A2(dbiEvent), .Z(n129));
Q_AN02 U523 ( .A0(n128), .A1(n122), .Z(callEmu));
Q_XOR2 U524 ( .A0(callEmuR), .A1(sendPO), .Z(n128));
Q_AN02 U525 ( .A0(sdlEnable), .A1(sdlStop), .Z(n127));
Q_AN02 U526 ( .A0(stop4), .A1(tbcEnable), .Z(n126));
Q_AN02 U527 ( .A0(stop2), .A1(tbcEnable), .Z(n125));
Q_AN02 U528 ( .A0(stop1), .A1(tbcEnable), .Z(n124));
Q_AN03 U529 ( .A0(n123), .A1(APPLY_PI), .A2(n122), .Z(dbiEvent));
Q_INV U530 ( .A(applyPiR), .Z(n123));
Q_INV U531 ( .A(hotSwapOnPI), .Z(n122));
Q_LDP0 \simTime_REG[0] ( .G(callEmu), .D(evalStepPI[0]), .Q(simTime[0]), .QN( ));
Q_LDP0 \simTime_REG[1] ( .G(callEmu), .D(evalStepPI[1]), .Q(simTime[1]), .QN( ));
Q_LDP0 \simTime_REG[2] ( .G(callEmu), .D(evalStepPI[2]), .Q(simTime[2]), .QN( ));
Q_LDP0 \simTime_REG[3] ( .G(callEmu), .D(evalStepPI[3]), .Q(simTime[3]), .QN( ));
Q_LDP0 \simTime_REG[4] ( .G(callEmu), .D(evalStepPI[4]), .Q(simTime[4]), .QN( ));
Q_LDP0 \simTime_REG[5] ( .G(callEmu), .D(evalStepPI[5]), .Q(simTime[5]), .QN( ));
Q_LDP0 \simTime_REG[6] ( .G(callEmu), .D(evalStepPI[6]), .Q(simTime[6]), .QN( ));
Q_LDP0 \simTime_REG[7] ( .G(callEmu), .D(evalStepPI[7]), .Q(simTime[7]), .QN( ));
Q_LDP0 \simTime_REG[8] ( .G(callEmu), .D(evalStepPI[8]), .Q(simTime[8]), .QN( ));
Q_LDP0 \simTime_REG[9] ( .G(callEmu), .D(evalStepPI[9]), .Q(simTime[9]), .QN( ));
Q_LDP0 \simTime_REG[10] ( .G(callEmu), .D(evalStepPI[10]), .Q(simTime[10]), .QN( ));
Q_LDP0 \simTime_REG[11] ( .G(callEmu), .D(evalStepPI[11]), .Q(simTime[11]), .QN( ));
Q_LDP0 \simTime_REG[12] ( .G(callEmu), .D(evalStepPI[12]), .Q(simTime[12]), .QN( ));
Q_LDP0 \simTime_REG[13] ( .G(callEmu), .D(evalStepPI[13]), .Q(simTime[13]), .QN( ));
Q_LDP0 \simTime_REG[14] ( .G(callEmu), .D(evalStepPI[14]), .Q(simTime[14]), .QN( ));
Q_LDP0 \simTime_REG[15] ( .G(callEmu), .D(evalStepPI[15]), .Q(simTime[15]), .QN( ));
Q_LDP0 \simTime_REG[16] ( .G(callEmu), .D(evalStepPI[16]), .Q(simTime[16]), .QN( ));
Q_LDP0 \simTime_REG[17] ( .G(callEmu), .D(evalStepPI[17]), .Q(simTime[17]), .QN( ));
Q_LDP0 \simTime_REG[18] ( .G(callEmu), .D(evalStepPI[18]), .Q(simTime[18]), .QN( ));
Q_LDP0 \simTime_REG[19] ( .G(callEmu), .D(evalStepPI[19]), .Q(simTime[19]), .QN( ));
Q_LDP0 \simTime_REG[20] ( .G(callEmu), .D(evalStepPI[20]), .Q(simTime[20]), .QN( ));
Q_LDP0 \simTime_REG[21] ( .G(callEmu), .D(evalStepPI[21]), .Q(simTime[21]), .QN( ));
Q_LDP0 \simTime_REG[22] ( .G(callEmu), .D(evalStepPI[22]), .Q(simTime[22]), .QN( ));
Q_LDP0 \simTime_REG[23] ( .G(callEmu), .D(evalStepPI[23]), .Q(simTime[23]), .QN( ));
Q_LDP0 \simTime_REG[24] ( .G(callEmu), .D(evalStepPI[24]), .Q(simTime[24]), .QN( ));
Q_LDP0 \simTime_REG[25] ( .G(callEmu), .D(evalStepPI[25]), .Q(simTime[25]), .QN( ));
Q_LDP0 \simTime_REG[26] ( .G(callEmu), .D(evalStepPI[26]), .Q(simTime[26]), .QN( ));
Q_LDP0 \simTime_REG[27] ( .G(callEmu), .D(evalStepPI[27]), .Q(simTime[27]), .QN( ));
Q_LDP0 \simTime_REG[28] ( .G(callEmu), .D(evalStepPI[28]), .Q(simTime[28]), .QN( ));
Q_LDP0 \simTime_REG[29] ( .G(callEmu), .D(evalStepPI[29]), .Q(simTime[29]), .QN( ));
Q_LDP0 \simTime_REG[30] ( .G(callEmu), .D(evalStepPI[30]), .Q(simTime[30]), .QN( ));
Q_LDP0 \simTime_REG[31] ( .G(callEmu), .D(evalStepPI[31]), .Q(simTime[31]), .QN( ));
Q_LDP0 \simTime_REG[32] ( .G(callEmu), .D(evalStepPI[32]), .Q(simTime[32]), .QN( ));
Q_LDP0 \simTime_REG[33] ( .G(callEmu), .D(evalStepPI[33]), .Q(simTime[33]), .QN( ));
Q_LDP0 \simTime_REG[34] ( .G(callEmu), .D(evalStepPI[34]), .Q(simTime[34]), .QN( ));
Q_LDP0 \simTime_REG[35] ( .G(callEmu), .D(evalStepPI[35]), .Q(simTime[35]), .QN( ));
Q_LDP0 \simTime_REG[36] ( .G(callEmu), .D(evalStepPI[36]), .Q(simTime[36]), .QN( ));
Q_LDP0 \simTime_REG[37] ( .G(callEmu), .D(evalStepPI[37]), .Q(simTime[37]), .QN( ));
Q_LDP0 \simTime_REG[38] ( .G(callEmu), .D(evalStepPI[38]), .Q(simTime[38]), .QN( ));
Q_LDP0 \simTime_REG[39] ( .G(callEmu), .D(evalStepPI[39]), .Q(simTime[39]), .QN( ));
Q_LDP0 \simTime_REG[40] ( .G(callEmu), .D(evalStepPI[40]), .Q(simTime[40]), .QN( ));
Q_LDP0 \simTime_REG[41] ( .G(callEmu), .D(evalStepPI[41]), .Q(simTime[41]), .QN( ));
Q_LDP0 \simTime_REG[42] ( .G(callEmu), .D(evalStepPI[42]), .Q(simTime[42]), .QN( ));
Q_LDP0 \simTime_REG[43] ( .G(callEmu), .D(evalStepPI[43]), .Q(simTime[43]), .QN( ));
Q_LDP0 \simTime_REG[44] ( .G(callEmu), .D(evalStepPI[44]), .Q(simTime[44]), .QN( ));
Q_LDP0 \simTime_REG[45] ( .G(callEmu), .D(evalStepPI[45]), .Q(simTime[45]), .QN( ));
Q_LDP0 \simTime_REG[46] ( .G(callEmu), .D(evalStepPI[46]), .Q(simTime[46]), .QN( ));
Q_LDP0 \simTime_REG[47] ( .G(callEmu), .D(evalStepPI[47]), .Q(simTime[47]), .QN( ));
Q_LDP0 \simTime_REG[48] ( .G(callEmu), .D(evalStepPI[48]), .Q(simTime[48]), .QN( ));
Q_LDP0 \simTime_REG[49] ( .G(callEmu), .D(evalStepPI[49]), .Q(simTime[49]), .QN( ));
Q_LDP0 \simTime_REG[50] ( .G(callEmu), .D(evalStepPI[50]), .Q(simTime[50]), .QN( ));
Q_LDP0 \simTime_REG[51] ( .G(callEmu), .D(evalStepPI[51]), .Q(simTime[51]), .QN( ));
Q_LDP0 \simTime_REG[52] ( .G(callEmu), .D(evalStepPI[52]), .Q(simTime[52]), .QN( ));
Q_LDP0 \simTime_REG[53] ( .G(callEmu), .D(evalStepPI[53]), .Q(simTime[53]), .QN( ));
Q_LDP0 \simTime_REG[54] ( .G(callEmu), .D(evalStepPI[54]), .Q(simTime[54]), .QN( ));
Q_LDP0 \simTime_REG[55] ( .G(callEmu), .D(evalStepPI[55]), .Q(simTime[55]), .QN( ));
Q_LDP0 \simTime_REG[56] ( .G(callEmu), .D(evalStepPI[56]), .Q(simTime[56]), .QN( ));
Q_LDP0 \simTime_REG[57] ( .G(callEmu), .D(evalStepPI[57]), .Q(simTime[57]), .QN( ));
Q_LDP0 \simTime_REG[58] ( .G(callEmu), .D(evalStepPI[58]), .Q(simTime[58]), .QN( ));
Q_LDP0 \simTime_REG[59] ( .G(callEmu), .D(evalStepPI[59]), .Q(simTime[59]), .QN( ));
Q_LDP0 \simTime_REG[60] ( .G(callEmu), .D(evalStepPI[60]), .Q(simTime[60]), .QN( ));
Q_LDP0 \simTime_REG[61] ( .G(callEmu), .D(evalStepPI[61]), .Q(simTime[61]), .QN( ));
Q_LDP0 \simTime_REG[62] ( .G(callEmu), .D(evalStepPI[62]), .Q(simTime[62]), .QN( ));
Q_LDP0 \simTime_REG[63] ( .G(callEmu), .D(evalStepPI[63]), .Q(simTime[63]), .QN( ));
Q_XNR2 U596 ( .A0(ckgHoldPI), .A1(eClkR), .Z(eClkv));
Q_OR03 U597 ( .A0(poDelay[7]), .A1(poDelay[6]), .A2(poDelay[5]), .Z(n116));
Q_OR03 U598 ( .A0(poDelay[4]), .A1(poDelay[3]), .A2(poDelay[2]), .Z(n117));
Q_OR03 U599 ( .A0(poDelay[1]), .A1(poDelay[0]), .A2(n116), .Z(n118));
Q_OR02 U600 ( .A0(n117), .A1(n118), .Z(poBusy));
Q_OR02 U601 ( .A0(lbrOn), .A1(hotSwapOnPI), .Z(lbrOnAll));
Q_NR03 U602 ( .A0(callEmu), .A1(dbiEvent), .A2(poBusy), .Z(intr));
Q_RDN U603 ( .Z(stop1));
Q_RDN U604 ( .Z(stop2));
Q_RDN U605 ( .Z(stop4));
Q_RDN U606 ( .Z(asyncCall));
Q_RDN U607 ( .Z(isfWait));
Q_RDN U608 ( .Z(osfWait));
Q_RDN U609 ( .Z(bWait));
Q_BUF U610 ( .A(_ET3_COMPILER_RESERVED_NAME_DBI_APPLY_), .Z(APPLY_PI));
Q_BUF U611 ( .A(lbrOnAll), .Z(_ET3_COMPILER_RESERVED_NAME_LBRKER_ON_));
Q_PULSE U612 ( .A(sendPO), .Z(rClk));
Q_PULSE U613 ( .A(eClkv), .Z(eClk));
ixc_assign intrBuf ( _ET3_COMPILER_RESERVED_NAME_ORION_INTERRUPT_, intr);
Q_RBUFZN  dum1 ( dummyW, n119, n120);
Q_RBUFZP  dum2 ( dummyW, n121, n1);
Q_INV U617 ( .A(remStepPO[63]), .Z(n2));
Q_FDP4EP \eCount_REG[63] ( .CK(rClk), .CE(n134), .R(n115), .D(n2), .Q(eCount[63]));
`ifdef CBV
reg [31:0] _zzcmds [0:15];
initial begin: U619
  integer i;
  for (i=0; i<=15; i=i+1) _zzcmds[i] =
`ifdef CBV_MEM_INIT1
  {32{1'b1}};
`else
  32'b0;
`endif
end
reg [31:0] n520;
buf(memWriteCmd, n520[0]);
always @(n115)
#0 begin
n520 = _zzcmds[{n115, n115, n115, n115}];
end
`else
MPR16X32 _zzcmds ( .A3(n115), .A2(n115), .A1(n115), .A0(n115), .SYNC_IN(n115), .DO31( ),
 .DO30( ), .DO29( ), .DO28( ), .DO27( ), .DO26( ), .DO25( ), .DO24( ), .DO23( ),
 .DO22( ), .DO21( ), .DO20( ), .DO19( ), .DO18( ), .DO17( ), .DO16( ), .DO15( ),
 .DO14( ), .DO13( ), .DO12( ), .DO11( ), .DO10( ), .DO9( ), .DO8( ), .DO7( ),
 .DO6( ), .DO5( ), .DO4( ), .DO3( ), .DO2( ), .DO1( ), .DO0(memWriteCmd), .SYNC_OUT( ));
// pragma CVASTRPROP INSTANCE "_zzcmds" HDL_MEMORY_DECL "1 31 0 0 15"
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "_zzcmds 1 31 0 0 15"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW16X32_MPR16X32
`else
module MPW16X32( A3, A2, A1, A0, DI31, DI30, DI29,
 DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21,
 DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5,
 DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A3, A2, A1, A0, DI31, DI30, DI29, DI28,
 DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18,
 DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8,
 DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR16X32_
`else
module MPR16X32( A3, A2, A1, A0, SYNC_IN, DO31, DO30,
 DO29, DO28, DO27, DO26, DO25, DO24, DO23, DO22,
 DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT);
input  A3, A2, A1, A0, SYNC_IN;
output  DO31, DO30, DO29, DO28, DO27, DO26, DO25, DO24,
 DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR16X32_
`endif
`define MPW16X32_MPR16X32
`endif
`endif
