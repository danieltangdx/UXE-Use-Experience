
module ASSERTION ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire FAILURE;
Q_ASSIGN U0 ( .B(xc_top.stop2), .A(FAILURE));
endmodule
