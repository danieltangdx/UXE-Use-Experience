architecture module of IXC_OSF is

begin
end module;
