architecture module of _ixc_isc is

begin
end module;
