architecture module of axis_busreg is
  component Q_BRP
    port(Z : out std_logic) ;
  end component ;

begin
  _UnNamed_Inst_10 : Q_BRP port map (z) ;
end module;
