// xc_work/v/6.sv
// /tools/cadence/UXE171_p98/tools.lnx86/etc/ixcom/IXCSF.sv:2
// NOTE: This file corresponds to a module in the Hardware/DUT partition
`timescale 1ps/100fs
module IXC_OSF_MB;
endmodule

