architecture module of ixc_ref is

begin
end module;
