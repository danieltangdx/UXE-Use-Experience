library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity _ixc_isc is
end _ixc_isc ;
