// xc_work/v/8.sv
// /tools/cadence/UXE171_p98/tools.lnx86/etc/ixcom/IXCSF.sv:444
// NOTE: This file corresponds to a module in the Hardware/DUT partition
`timescale 1ps/100fs
module IXC_OSF1;
endmodule

