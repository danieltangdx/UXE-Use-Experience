architecture module of IXC_OSF1 is

begin
end module;
