module counter_tb;
 counter dut();
endmodule

