architecture module of ixc_assign is

begin

  process --:o822
  (*)
  begin
    L <= R ;
  end process ;
end module;
