
module IXC_MC_IFIFO ( ackClkX, ackLenX);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output ackClkX;
output [17:0] ackLenX;
wire ackClk;
wire ackClkN;
wire [17:0] ackLen;
wire [15:0] tId;
wire [511:0] iData;
wire [16:0] wptr;
wire [16:0] wptrN;
wire [16:0] xptr;
wire [16:0] xptrN;
wire [255:0] afifoXdata;
wire [255:0] afifoXdataFinal;
wire [16:0] rptr;
wire [16:0] rptrN;
wire [14:0] afifoRaddr0;
wire [14:0] afifoRaddr1;
wire [14:0] afifoRaddr2;
wire [767:0] afifoRdata;
wire [17:0] rdDelta;
wire [63:0] afifoRdCnt;
wire [3:0] markBits;
wire [3:0] markBitsN;
wire [3:0] newMarkBits;
wire [3:0] newMarkBitsD;
wire [3:0] dataBits;
wire [23:0] offset;
wire [23:0] offsetN;
wire moveForward;
wire moveForwardN;
wire active;
wire activeD;
wire [63:0] xval;
wire nps;
wire eob;
wire SFIFOLock;
wire [31:0] i;
wire [63:0] head;
wire [63:0] xhead;
wire [63:0] vhead;
wire [15:0] pktl;
wire [15:0] pktlN;
wire [15:0] vlen;
wire [15:0] vlenN;
wire rstDone;
wire rstDoneD;
wire rstDoneD2;
wire rstDoneD3;
wire rstDoneD4;
wire [11:0] odly;
wire [11:0] odlyN;
wire vmode;
wire [575:0] tmpData;
wire oSt;
wire [63:0] oMark;
wire [511:0] oData;
wire [511:0] oDataD;
wire [511:0] oDataD2;
wire oDataEn;
wire oDataEnD;
wire oDataEnD2;
wire [3:0] oDataLen;
wire [3:0] oDataLenD;
wire [3:0] oDataLenD2;
wire [767:0] bfifoData;
wire [3:0] bFill;
wire [14:0] bfifoAddr0;
wire [15:0] bfifoAddr1;
wire [15:0] bfifoAddr2;
wire [14:0] bfifoWptr;
wire [7:0] shiftCount;
wire [767:0] shiftedOData;
Q_NOT_TOUCH _zzqnthw ( .sig(n1));
endmodule
