ARCHITECTURE module OF ixc_assign_32 IS

BEGIN

  PROCESS --:o822
  (*)
  BEGIN
    L <= R ;
  END PROCESS ;
END module;