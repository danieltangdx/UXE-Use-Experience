architecture module of ixc_asgn_cov_rst_pulse is
  signal DUMMY0 : std_logic ;

begin
  rstsig <= DUMMY0 ;
end module;
