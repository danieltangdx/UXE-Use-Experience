architecture module of ixc_frequency is
  -- quickturn CVASTRPROP MODULE HDLICE IXCOM_FREQUENCY_CELL "1"

begin
end module;
