
module counter ( clk, out);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
output [31:0] out;
wire [31:0] counter;
supply0 n62;
ixc_assign_32 _zz_strnp_1 ( out[31:0], counter[31:0]);
Q_FDP0 \counter_REG[0] ( .CK(clk), .D(n61), .Q(counter[0]), .QN(n61));
Q_FDP0 \counter_REG[1] ( .CK(clk), .D(n60), .Q(counter[1]), .QN( ));
Q_FDP0 \counter_REG[2] ( .CK(clk), .D(n58), .Q(counter[2]), .QN( ));
Q_FDP0 \counter_REG[3] ( .CK(clk), .D(n56), .Q(counter[3]), .QN( ));
Q_FDP0 \counter_REG[4] ( .CK(clk), .D(n54), .Q(counter[4]), .QN( ));
Q_FDP0 \counter_REG[5] ( .CK(clk), .D(n52), .Q(counter[5]), .QN( ));
Q_FDP0 \counter_REG[6] ( .CK(clk), .D(n50), .Q(counter[6]), .QN( ));
Q_FDP0 \counter_REG[7] ( .CK(clk), .D(n48), .Q(counter[7]), .QN( ));
Q_FDP0 \counter_REG[8] ( .CK(clk), .D(n46), .Q(counter[8]), .QN( ));
Q_FDP0 \counter_REG[9] ( .CK(clk), .D(n44), .Q(counter[9]), .QN( ));
Q_FDP0 \counter_REG[10] ( .CK(clk), .D(n42), .Q(counter[10]), .QN( ));
Q_FDP0 \counter_REG[11] ( .CK(clk), .D(n40), .Q(counter[11]), .QN( ));
Q_FDP0 \counter_REG[12] ( .CK(clk), .D(n38), .Q(counter[12]), .QN( ));
Q_FDP0 \counter_REG[13] ( .CK(clk), .D(n36), .Q(counter[13]), .QN( ));
Q_FDP0 \counter_REG[14] ( .CK(clk), .D(n34), .Q(counter[14]), .QN( ));
Q_FDP0 \counter_REG[15] ( .CK(clk), .D(n32), .Q(counter[15]), .QN( ));
Q_FDP0 \counter_REG[16] ( .CK(clk), .D(n30), .Q(counter[16]), .QN( ));
Q_FDP0 \counter_REG[17] ( .CK(clk), .D(n28), .Q(counter[17]), .QN( ));
Q_FDP0 \counter_REG[18] ( .CK(clk), .D(n26), .Q(counter[18]), .QN( ));
Q_FDP0 \counter_REG[19] ( .CK(clk), .D(n24), .Q(counter[19]), .QN( ));
Q_FDP0 \counter_REG[20] ( .CK(clk), .D(n22), .Q(counter[20]), .QN( ));
Q_FDP0 \counter_REG[21] ( .CK(clk), .D(n20), .Q(counter[21]), .QN( ));
Q_FDP0 \counter_REG[22] ( .CK(clk), .D(n18), .Q(counter[22]), .QN( ));
Q_FDP0 \counter_REG[23] ( .CK(clk), .D(n16), .Q(counter[23]), .QN( ));
Q_FDP0 \counter_REG[24] ( .CK(clk), .D(n14), .Q(counter[24]), .QN( ));
Q_FDP0 \counter_REG[25] ( .CK(clk), .D(n12), .Q(counter[25]), .QN( ));
Q_FDP0 \counter_REG[26] ( .CK(clk), .D(n10), .Q(counter[26]), .QN( ));
Q_FDP0 \counter_REG[27] ( .CK(clk), .D(n8), .Q(counter[27]), .QN( ));
Q_FDP0 \counter_REG[28] ( .CK(clk), .D(n6), .Q(counter[28]), .QN( ));
Q_FDP0 \counter_REG[29] ( .CK(clk), .D(n4), .Q(counter[29]), .QN( ));
Q_FDP0 \counter_REG[30] ( .CK(clk), .D(n2), .Q(counter[30]), .QN( ));
Q_AD01HF U32 ( .A0(counter[30]), .B0(n3), .S(n2), .CO(n1));
Q_AD01HF U33 ( .A0(counter[29]), .B0(n5), .S(n4), .CO(n3));
Q_AD01HF U34 ( .A0(counter[28]), .B0(n7), .S(n6), .CO(n5));
Q_AD01HF U35 ( .A0(counter[27]), .B0(n9), .S(n8), .CO(n7));
Q_AD01HF U36 ( .A0(counter[26]), .B0(n11), .S(n10), .CO(n9));
Q_AD01HF U37 ( .A0(counter[25]), .B0(n13), .S(n12), .CO(n11));
Q_AD01HF U38 ( .A0(counter[24]), .B0(n15), .S(n14), .CO(n13));
Q_AD01HF U39 ( .A0(counter[23]), .B0(n17), .S(n16), .CO(n15));
Q_AD01HF U40 ( .A0(counter[22]), .B0(n19), .S(n18), .CO(n17));
Q_AD01HF U41 ( .A0(counter[21]), .B0(n21), .S(n20), .CO(n19));
Q_AD01HF U42 ( .A0(counter[20]), .B0(n23), .S(n22), .CO(n21));
Q_AD01HF U43 ( .A0(counter[19]), .B0(n25), .S(n24), .CO(n23));
Q_AD01HF U44 ( .A0(counter[18]), .B0(n27), .S(n26), .CO(n25));
Q_AD01HF U45 ( .A0(counter[17]), .B0(n29), .S(n28), .CO(n27));
Q_AD01HF U46 ( .A0(counter[16]), .B0(n31), .S(n30), .CO(n29));
Q_AD01HF U47 ( .A0(counter[15]), .B0(n33), .S(n32), .CO(n31));
Q_AD01HF U48 ( .A0(counter[14]), .B0(n35), .S(n34), .CO(n33));
Q_AD01HF U49 ( .A0(counter[13]), .B0(n37), .S(n36), .CO(n35));
Q_AD01HF U50 ( .A0(counter[12]), .B0(n39), .S(n38), .CO(n37));
Q_AD01HF U51 ( .A0(counter[11]), .B0(n41), .S(n40), .CO(n39));
Q_AD01HF U52 ( .A0(counter[10]), .B0(n43), .S(n42), .CO(n41));
Q_AD01HF U53 ( .A0(counter[9]), .B0(n45), .S(n44), .CO(n43));
Q_AD01HF U54 ( .A0(counter[8]), .B0(n47), .S(n46), .CO(n45));
Q_AD01HF U55 ( .A0(counter[7]), .B0(n49), .S(n48), .CO(n47));
Q_AD01HF U56 ( .A0(counter[6]), .B0(n51), .S(n50), .CO(n49));
Q_AD01HF U57 ( .A0(counter[5]), .B0(n53), .S(n52), .CO(n51));
Q_AD01HF U58 ( .A0(counter[4]), .B0(n55), .S(n54), .CO(n53));
Q_AD01HF U59 ( .A0(counter[3]), .B0(n57), .S(n56), .CO(n55));
Q_AD01HF U60 ( .A0(counter[2]), .B0(n59), .S(n58), .CO(n57));
Q_AD01HF U61 ( .A0(counter[1]), .B0(counter[0]), .S(n60), .CO(n59));
Q_INV U62 ( .A(counter[31]), .Z(n63));
Q_FDP4EP \counter_REG[31] ( .CK(clk), .CE(n1), .R(n62), .D(n63), .Q(counter[31]));
endmodule
