architecture module of IXC_OSF_MB is

begin
end module;
